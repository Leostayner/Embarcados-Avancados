-- nioshello_ps2_0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity nioshello_ps2_0 is
	generic (
		LEN : natural := 4
	);
	port (
		clk           : in    std_logic                     := '0';             --          clock.clk
		reset         : in    std_logic                     := '0';             --          reset.reset
		avs_address   : in    std_logic_vector(3 downto 0)  := (others => '0'); -- avalon_slave_0.address
		avs_read      : in    std_logic                     := '0';             --               .read
		avs_readdata  : out   std_logic_vector(31 downto 0);                    --               .readdata
		avs_write     : in    std_logic                     := '0';             --               .write
		avs_writedata : in    std_logic_vector(31 downto 0) := (others => '0'); --               .writedata
		PS2_CLK       : inout std_logic                     := '0';             --            clk.export
		PS2_DAT       : inout std_logic                     := '0'              --            dat.export
	);
end entity nioshello_ps2_0;

architecture rtl of nioshello_ps2_0 is
	component peripheral_LED is
		generic (
			LEN : natural := 4
		);
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			reset         : in    std_logic                     := 'X';             -- reset
			avs_address   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			avs_read      : in    std_logic                     := 'X';             -- read
			avs_readdata  : out   std_logic_vector(31 downto 0);                    -- readdata
			avs_write     : in    std_logic                     := 'X';             -- write
			avs_writedata : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			PS2_CLK       : inout std_logic                     := 'X';             -- export
			PS2_DAT       : inout std_logic                     := 'X'              -- export
		);
	end component peripheral_LED;

begin

	len_check : if LEN /= 4 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	ps2_0 : component peripheral_LED
		generic map (
			LEN => 4
		)
		port map (
			clk           => clk,           --          clock.clk
			reset         => reset,         --          reset.reset
			avs_address   => avs_address,   -- avalon_slave_0.address
			avs_read      => avs_read,      --               .read
			avs_readdata  => avs_readdata,  --               .readdata
			avs_write     => avs_write,     --               .write
			avs_writedata => avs_writedata, --               .writedata
			PS2_CLK       => PS2_CLK,       --            clk.export
			PS2_DAT       => PS2_DAT        --            dat.export
		);

end architecture rtl; -- of nioshello_ps2_0
